library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity RSA is
    port(

    );
end RSA;

architecture internal of RSA is

begin

end architecture;